module or_gate_bit (input a, b,
               output cout);
  assign cout = a | b;
endmodule
