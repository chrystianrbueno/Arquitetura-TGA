module and_gate (a, b, cout);
 input a, b;
 output cout;
 assign cout = a & b;
endmodule